.title KiCad schematic
.include "models/XLamp-XBD-Spice.txt"
V1 /IN 0 {VIN}
D1 /IN /BRANCH01 XB-DWHT
D2 /IN /BRANCH01 XB-DWHT
D4 /BRANCH01 /BRANCH02 XB-DWHT
D5 /BRANCH01 /BRANCH02 XB-DWHT
D7 /BRANCH02 /BRANCH03 XB-DWHT
D8 /BRANCH02 /BRANCH03 XB-DWHT
D10 /BRANCH03 /BRANCH04 XB-DWHT
D11 /BRANCH03 /BRANCH04 XB-DWHT
D13 /BRANCH04 /BRANCH05 XB-DWHT
D14 /BRANCH04 /BRANCH05 XB-DWHT
D16 /BRANCH05 /BRANCH06 XB-DWHT
D17 /BRANCH05 /BRANCH06 XB-DWHT
D3 /IN /BRANCH01 XB-DWHT
D6 /BRANCH01 /BRANCH02 XB-DWHT
D9 /BRANCH02 /BRANCH03 XB-DWHT
D12 /BRANCH03 /BRANCH04 XB-DWHT
D15 /BRANCH04 /BRANCH05 XB-DWHT
D18 /BRANCH05 /BRANCH06 XB-DWHT
D19 /BRANCH06 0 XB-DWHT
D20 /BRANCH06 0 XB-DWHT
D21 /BRANCH06 0 XB-DWHT
.end
